** sch_path: /home/shahid/Sky130Projects/inv/Xschem/inv_tb.sch
**.subckt inv_tb
x1 VSS VDD OUT IN inv
V1 VSS GND 0
V2 VDD VSS 1.8
V3 IN VSS pulse(0 1.8 0 100p 100p 100n 200n)
C1 OUT VSS 20f m=1
*  CORNER -  corner  IS MISSING !!!!
**** begin user architecture code

* this option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1
.option savecurrents
.control
save all

dc v3 0 1.8 0.025
plot v(IN) v(OUT)

tran 10p 1u
plot v(IN) v(OUT)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/shahid/Sky130Projects/inv/Xschem/inv.sym
** sch_path: /home/shahid/Sky130Projects/inv/Xschem/inv.sch
.subckt inv VSS VDD OUT IN
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
*  M1 -  nfet_01v8  IS MISSING !!!!
*  M2 -  pfet_01v8  IS MISSING !!!!
.ends

.GLOBAL GND
.end
