* NGSPICE file created from INV_MAG_flat.ext - technology: sky130A

.subckt inv_pex VSS VDD OUT IN
X0 OUT.t3 IN.t0 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 OUT.t2 IN.t1 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2 OUT.t0 IN.t2 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 OUT.t1 IN.t3 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
R0 IN.n0 IN.t0 468.464
R1 IN.n2 IN.t1 308.428
R2 IN.n1 IN.t3 284.38
R3 IN.n0 IN.t2 249.034
R4 IN.n2 IN.n1 83.9618
R5 IN IN.n2 44.0365
R6 IN.n1 IN.n0 14.4605
R7 VDD.t0 VDD.t2 479.399
R8 VDD.n0 VDD.t4 475
R9 VDD.n4 VDD.t3 128.312
R10 VDD.n3 VDD.t5 120.135
R11 VDD.n4 VDD.t1 89.5567
R12 VDD.n2 VDD.n1 43.3338
R13 VDD VDD.n3 4.62272
R14 VDD.n0 VDD.t0 4.39865
R15 VDD VDD.n4 3.55606
R16 VDD.n3 VDD.n2 0.000536524
R17 VDD.n2 VDD.n0 0.000536524
R18 OUT.n0 OUT.t2 29.5446
R19 OUT.n1 OUT.t3 29.0103
R20 OUT.n0 OUT.t1 29.0103
R21 OUT.n0 OUT.t0 17.7528
R22 OUT.n1 OUT.n0 0.534814
R23 OUT OUT.n1 0.145108
R24 VSS.n1 VSS.t0 1352.29
R25 VSS VSS.t1 87.1655
R26 VSS.n1 VSS.n0 1.36618
R27 VSS VSS.n1 0.356217
C0 VDD OUT 0.864f
C1 OUT IN 0.143f
C2 VDD IN 0.342f
.ends

