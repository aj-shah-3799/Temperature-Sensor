** sch_path: /home/shahid/Sky130Projects/inv/Xschem/inv _pex_tb.sch
**.subckt inv _pex_tb
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 1.8
.save i(v2)
V3 IN VSS pulse(0 1.8 0 100p 100p 100n 200n)
.save i(v3)
C1 OUT VSS 20f m=1
x1 VSS VDD OUT IN inv_pex
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


* this option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1
.option savecurrents
.include pex_INV_MAG.spice
.control
save all

dc v3 0 1.8 0.025
plot v(IN) v(OUT)

tran 10p 1u
plot v(IN) v(OUT)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
